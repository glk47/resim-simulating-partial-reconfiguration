------------------------------------------------------------------------------
-- THIS FILE IS EMPTY BUT CAN NOT BE DELETED
------------------------------------------------------------------------------
